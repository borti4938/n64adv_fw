//////////////////////////////////////////////////////////////////////////////////
//
// This file is part of the N64 RGB/YPbPr DAC project.
//
// Copyright (C) 2015-2022 by Peter Bartmann <borti4938@gmail.com>
//
// N64 RGB/YPbPr DAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//////////////////////////////////////////////////////////////////////////////////
//
// Company:  Circuit-Board.de
// Engineer: borti4938
//
// Module Name:    font_rom
// Project Name:   N64 Advanced RGB/YPbPr DAC Mod
// Target Devices: Max10, Cyclone IV and Cyclone 10 LP devices
// Tool versions:  Altera Quartus Prime
// Description:    simple line-multiplying
//
// Features: ip independent implementation of font rom
//
// This file is auto generated by script/font2rom.m
//
//////////////////////////////////////////////////////////////////////////////////


module font_rom(
  CLK,
  nRST,
  char_addr,
  char_line,
  rden,
  rddata
);

input       CLK;
input       nRST;
input [6:0] char_addr;
input [3:0] char_line;
input       rden;

output reg [7:0] rddata = 8'h0;


reg [10:0] addr_r = 11'h00;
reg        rden_r =  1'b0;

reg [7:0] font_mem[0:1535];
initial begin
  font_mem[0000] = 000;
  font_mem[0001] = 000;
  font_mem[0002] = 000;
  font_mem[0003] = 000;
  font_mem[0004] = 000;
  font_mem[0005] = 000;
  font_mem[0006] = 000;
  font_mem[0007] = 000;
  font_mem[0008] = 000;
  font_mem[0009] = 000;
  font_mem[0010] = 000;
  font_mem[0011] = 000;
  font_mem[0012] = 000;
  font_mem[0013] = 000;
  font_mem[0014] = 000;
  font_mem[0015] = 000;
  font_mem[0016] = 000;
  font_mem[0017] = 000;
  font_mem[0018] = 000;
  font_mem[0019] = 000;
  font_mem[0020] = 000;
  font_mem[0021] = 000;
  font_mem[0022] = 000;
  font_mem[0023] = 000;
  font_mem[0024] = 000;
  font_mem[0025] = 000;
  font_mem[0026] = 000;
  font_mem[0027] = 000;
  font_mem[0028] = 000;
  font_mem[0029] = 000;
  font_mem[0030] = 000;
  font_mem[0031] = 000;
  font_mem[0032] = 000;
  font_mem[0033] = 000;
  font_mem[0034] = 000;
  font_mem[0035] = 000;
  font_mem[0036] = 012;
  font_mem[0037] = 000;
  font_mem[0038] = 000;
  font_mem[0039] = 000;
  font_mem[0040] = 000;
  font_mem[0041] = 000;
  font_mem[0042] = 000;
  font_mem[0043] = 000;
  font_mem[0044] = 000;
  font_mem[0045] = 000;
  font_mem[0046] = 000;
  font_mem[0047] = 000;
  font_mem[0048] = 000;
  font_mem[0049] = 000;
  font_mem[0050] = 000;
  font_mem[0051] = 000;
  font_mem[0052] = 000;
  font_mem[0053] = 000;
  font_mem[0054] = 000;
  font_mem[0055] = 000;
  font_mem[0056] = 000;
  font_mem[0057] = 000;
  font_mem[0058] = 000;
  font_mem[0059] = 000;
  font_mem[0060] = 000;
  font_mem[0061] = 000;
  font_mem[0062] = 000;
  font_mem[0063] = 000;
  font_mem[0064] = 000;
  font_mem[0065] = 000;
  font_mem[0066] = 000;
  font_mem[0067] = 000;
  font_mem[0068] = 000;
  font_mem[0069] = 000;
  font_mem[0070] = 000;
  font_mem[0071] = 000;
  font_mem[0072] = 000;
  font_mem[0073] = 000;
  font_mem[0074] = 000;
  font_mem[0075] = 000;
  font_mem[0076] = 000;
  font_mem[0077] = 000;
  font_mem[0078] = 000;
  font_mem[0079] = 000;
  font_mem[0080] = 000;
  font_mem[0081] = 000;
  font_mem[0082] = 000;
  font_mem[0083] = 000;
  font_mem[0084] = 000;
  font_mem[0085] = 000;
  font_mem[0086] = 000;
  font_mem[0087] = 000;
  font_mem[0088] = 000;
  font_mem[0089] = 000;
  font_mem[0090] = 000;
  font_mem[0091] = 000;
  font_mem[0092] = 000;
  font_mem[0093] = 000;
  font_mem[0094] = 008;
  font_mem[0095] = 000;
  font_mem[0096] = 012;
  font_mem[0097] = 000;
  font_mem[0098] = 000;
  font_mem[0099] = 000;
  font_mem[0100] = 000;
  font_mem[0101] = 000;
  font_mem[0102] = 000;
  font_mem[0103] = 000;
  font_mem[0104] = 000;
  font_mem[0105] = 000;
  font_mem[0106] = 000;
  font_mem[0107] = 000;
  font_mem[0108] = 000;
  font_mem[0109] = 000;
  font_mem[0110] = 000;
  font_mem[0111] = 000;
  font_mem[0112] = 000;
  font_mem[0113] = 000;
  font_mem[0114] = 000;
  font_mem[0115] = 000;
  font_mem[0116] = 000;
  font_mem[0117] = 000;
  font_mem[0118] = 000;
  font_mem[0119] = 000;
  font_mem[0120] = 000;
  font_mem[0121] = 000;
  font_mem[0122] = 000;
  font_mem[0123] = 000;
  font_mem[0124] = 000;
  font_mem[0125] = 000;
  font_mem[0126] = 000;
  font_mem[0127] = 000;
  font_mem[0128] = 000;
  font_mem[0129] = 000;
  font_mem[0130] = 126;
  font_mem[0131] = 000;
  font_mem[0132] = 008;
  font_mem[0133] = 024;
  font_mem[0134] = 024;
  font_mem[0135] = 000;
  font_mem[0136] = 000;
  font_mem[0137] = 028;
  font_mem[0138] = 028;
  font_mem[0139] = 124;
  font_mem[0140] = 060;
  font_mem[0141] = 000;
  font_mem[0142] = 254;
  font_mem[0143] = 000;
  font_mem[0144] = 064;
  font_mem[0145] = 001;
  font_mem[0146] = 024;
  font_mem[0147] = 102;
  font_mem[0148] = 254;
  font_mem[0149] = 126;
  font_mem[0150] = 000;
  font_mem[0151] = 024;
  font_mem[0152] = 024;
  font_mem[0153] = 024;
  font_mem[0154] = 000;
  font_mem[0155] = 000;
  font_mem[0156] = 000;
  font_mem[0157] = 000;
  font_mem[0158] = 000;
  font_mem[0159] = 000;
  font_mem[0160] = 000;
  font_mem[0161] = 012;
  font_mem[0162] = 102;
  font_mem[0163] = 054;
  font_mem[0164] = 012;
  font_mem[0165] = 000;
  font_mem[0166] = 014;
  font_mem[0167] = 012;
  font_mem[0168] = 048;
  font_mem[0169] = 006;
  font_mem[0170] = 000;
  font_mem[0171] = 000;
  font_mem[0172] = 000;
  font_mem[0173] = 000;
  font_mem[0174] = 000;
  font_mem[0175] = 000;
  font_mem[0176] = 062;
  font_mem[0177] = 008;
  font_mem[0178] = 030;
  font_mem[0179] = 030;
  font_mem[0180] = 048;
  font_mem[0181] = 063;
  font_mem[0182] = 028;
  font_mem[0183] = 127;
  font_mem[0184] = 030;
  font_mem[0185] = 030;
  font_mem[0186] = 000;
  font_mem[0187] = 000;
  font_mem[0188] = 048;
  font_mem[0189] = 000;
  font_mem[0190] = 006;
  font_mem[0191] = 030;
  font_mem[0192] = 062;
  font_mem[0193] = 012;
  font_mem[0194] = 063;
  font_mem[0195] = 060;
  font_mem[0196] = 031;
  font_mem[0197] = 127;
  font_mem[0198] = 127;
  font_mem[0199] = 060;
  font_mem[0200] = 051;
  font_mem[0201] = 030;
  font_mem[0202] = 120;
  font_mem[0203] = 103;
  font_mem[0204] = 015;
  font_mem[0205] = 099;
  font_mem[0206] = 099;
  font_mem[0207] = 028;
  font_mem[0208] = 063;
  font_mem[0209] = 028;
  font_mem[0210] = 063;
  font_mem[0211] = 030;
  font_mem[0212] = 063;
  font_mem[0213] = 051;
  font_mem[0214] = 051;
  font_mem[0215] = 099;
  font_mem[0216] = 051;
  font_mem[0217] = 051;
  font_mem[0218] = 127;
  font_mem[0219] = 060;
  font_mem[0220] = 000;
  font_mem[0221] = 060;
  font_mem[0222] = 028;
  font_mem[0223] = 000;
  font_mem[0224] = 012;
  font_mem[0225] = 000;
  font_mem[0226] = 007;
  font_mem[0227] = 000;
  font_mem[0228] = 056;
  font_mem[0229] = 000;
  font_mem[0230] = 028;
  font_mem[0231] = 000;
  font_mem[0232] = 007;
  font_mem[0233] = 024;
  font_mem[0234] = 048;
  font_mem[0235] = 007;
  font_mem[0236] = 030;
  font_mem[0237] = 000;
  font_mem[0238] = 000;
  font_mem[0239] = 000;
  font_mem[0240] = 000;
  font_mem[0241] = 000;
  font_mem[0242] = 000;
  font_mem[0243] = 000;
  font_mem[0244] = 000;
  font_mem[0245] = 000;
  font_mem[0246] = 000;
  font_mem[0247] = 000;
  font_mem[0248] = 000;
  font_mem[0249] = 000;
  font_mem[0250] = 000;
  font_mem[0251] = 056;
  font_mem[0252] = 024;
  font_mem[0253] = 007;
  font_mem[0254] = 206;
  font_mem[0255] = 000;
  font_mem[0256] = 000;
  font_mem[0257] = 000;
  font_mem[0258] = 195;
  font_mem[0259] = 034;
  font_mem[0260] = 028;
  font_mem[0261] = 060;
  font_mem[0262] = 060;
  font_mem[0263] = 255;
  font_mem[0264] = 255;
  font_mem[0265] = 034;
  font_mem[0266] = 034;
  font_mem[0267] = 112;
  font_mem[0268] = 102;
  font_mem[0269] = 000;
  font_mem[0270] = 198;
  font_mem[0271] = 024;
  font_mem[0272] = 096;
  font_mem[0273] = 003;
  font_mem[0274] = 060;
  font_mem[0275] = 102;
  font_mem[0276] = 219;
  font_mem[0277] = 198;
  font_mem[0278] = 000;
  font_mem[0279] = 060;
  font_mem[0280] = 060;
  font_mem[0281] = 024;
  font_mem[0282] = 000;
  font_mem[0283] = 000;
  font_mem[0284] = 000;
  font_mem[0285] = 000;
  font_mem[0286] = 008;
  font_mem[0287] = 127;
  font_mem[0288] = 000;
  font_mem[0289] = 030;
  font_mem[0290] = 102;
  font_mem[0291] = 054;
  font_mem[0292] = 062;
  font_mem[0293] = 000;
  font_mem[0294] = 027;
  font_mem[0295] = 012;
  font_mem[0296] = 024;
  font_mem[0297] = 012;
  font_mem[0298] = 000;
  font_mem[0299] = 000;
  font_mem[0300] = 000;
  font_mem[0301] = 000;
  font_mem[0302] = 000;
  font_mem[0303] = 064;
  font_mem[0304] = 099;
  font_mem[0305] = 012;
  font_mem[0306] = 051;
  font_mem[0307] = 051;
  font_mem[0308] = 056;
  font_mem[0309] = 003;
  font_mem[0310] = 006;
  font_mem[0311] = 099;
  font_mem[0312] = 051;
  font_mem[0313] = 051;
  font_mem[0314] = 000;
  font_mem[0315] = 000;
  font_mem[0316] = 024;
  font_mem[0317] = 000;
  font_mem[0318] = 012;
  font_mem[0319] = 051;
  font_mem[0320] = 099;
  font_mem[0321] = 030;
  font_mem[0322] = 102;
  font_mem[0323] = 102;
  font_mem[0324] = 054;
  font_mem[0325] = 070;
  font_mem[0326] = 102;
  font_mem[0327] = 102;
  font_mem[0328] = 051;
  font_mem[0329] = 012;
  font_mem[0330] = 048;
  font_mem[0331] = 102;
  font_mem[0332] = 006;
  font_mem[0333] = 119;
  font_mem[0334] = 099;
  font_mem[0335] = 054;
  font_mem[0336] = 102;
  font_mem[0337] = 054;
  font_mem[0338] = 102;
  font_mem[0339] = 051;
  font_mem[0340] = 045;
  font_mem[0341] = 051;
  font_mem[0342] = 051;
  font_mem[0343] = 099;
  font_mem[0344] = 051;
  font_mem[0345] = 051;
  font_mem[0346] = 115;
  font_mem[0347] = 012;
  font_mem[0348] = 001;
  font_mem[0349] = 048;
  font_mem[0350] = 054;
  font_mem[0351] = 000;
  font_mem[0352] = 024;
  font_mem[0353] = 000;
  font_mem[0354] = 006;
  font_mem[0355] = 000;
  font_mem[0356] = 048;
  font_mem[0357] = 000;
  font_mem[0358] = 054;
  font_mem[0359] = 000;
  font_mem[0360] = 006;
  font_mem[0361] = 024;
  font_mem[0362] = 048;
  font_mem[0363] = 006;
  font_mem[0364] = 024;
  font_mem[0365] = 000;
  font_mem[0366] = 000;
  font_mem[0367] = 000;
  font_mem[0368] = 000;
  font_mem[0369] = 000;
  font_mem[0370] = 000;
  font_mem[0371] = 000;
  font_mem[0372] = 004;
  font_mem[0373] = 000;
  font_mem[0374] = 000;
  font_mem[0375] = 000;
  font_mem[0376] = 000;
  font_mem[0377] = 000;
  font_mem[0378] = 000;
  font_mem[0379] = 012;
  font_mem[0380] = 024;
  font_mem[0381] = 012;
  font_mem[0382] = 091;
  font_mem[0383] = 000;
  font_mem[0384] = 000;
  font_mem[0385] = 000;
  font_mem[0386] = 129;
  font_mem[0387] = 119;
  font_mem[0388] = 062;
  font_mem[0389] = 060;
  font_mem[0390] = 126;
  font_mem[0391] = 000;
  font_mem[0392] = 000;
  font_mem[0393] = 093;
  font_mem[0394] = 093;
  font_mem[0395] = 092;
  font_mem[0396] = 102;
  font_mem[0397] = 099;
  font_mem[0398] = 254;
  font_mem[0399] = 219;
  font_mem[0400] = 112;
  font_mem[0401] = 007;
  font_mem[0402] = 126;
  font_mem[0403] = 102;
  font_mem[0404] = 219;
  font_mem[0405] = 012;
  font_mem[0406] = 000;
  font_mem[0407] = 126;
  font_mem[0408] = 126;
  font_mem[0409] = 024;
  font_mem[0410] = 012;
  font_mem[0411] = 024;
  font_mem[0412] = 000;
  font_mem[0413] = 036;
  font_mem[0414] = 008;
  font_mem[0415] = 127;
  font_mem[0416] = 000;
  font_mem[0417] = 030;
  font_mem[0418] = 102;
  font_mem[0419] = 127;
  font_mem[0420] = 003;
  font_mem[0421] = 035;
  font_mem[0422] = 027;
  font_mem[0423] = 012;
  font_mem[0424] = 012;
  font_mem[0425] = 024;
  font_mem[0426] = 102;
  font_mem[0427] = 024;
  font_mem[0428] = 000;
  font_mem[0429] = 000;
  font_mem[0430] = 000;
  font_mem[0431] = 096;
  font_mem[0432] = 115;
  font_mem[0433] = 015;
  font_mem[0434] = 051;
  font_mem[0435] = 048;
  font_mem[0436] = 060;
  font_mem[0437] = 003;
  font_mem[0438] = 003;
  font_mem[0439] = 099;
  font_mem[0440] = 051;
  font_mem[0441] = 051;
  font_mem[0442] = 028;
  font_mem[0443] = 028;
  font_mem[0444] = 012;
  font_mem[0445] = 000;
  font_mem[0446] = 024;
  font_mem[0447] = 048;
  font_mem[0448] = 099;
  font_mem[0449] = 051;
  font_mem[0450] = 102;
  font_mem[0451] = 099;
  font_mem[0452] = 102;
  font_mem[0453] = 006;
  font_mem[0454] = 070;
  font_mem[0455] = 099;
  font_mem[0456] = 051;
  font_mem[0457] = 012;
  font_mem[0458] = 048;
  font_mem[0459] = 054;
  font_mem[0460] = 006;
  font_mem[0461] = 127;
  font_mem[0462] = 103;
  font_mem[0463] = 099;
  font_mem[0464] = 102;
  font_mem[0465] = 099;
  font_mem[0466] = 102;
  font_mem[0467] = 051;
  font_mem[0468] = 012;
  font_mem[0469] = 051;
  font_mem[0470] = 051;
  font_mem[0471] = 099;
  font_mem[0472] = 051;
  font_mem[0473] = 051;
  font_mem[0474] = 025;
  font_mem[0475] = 012;
  font_mem[0476] = 003;
  font_mem[0477] = 048;
  font_mem[0478] = 099;
  font_mem[0479] = 000;
  font_mem[0480] = 000;
  font_mem[0481] = 000;
  font_mem[0482] = 006;
  font_mem[0483] = 000;
  font_mem[0484] = 048;
  font_mem[0485] = 000;
  font_mem[0486] = 006;
  font_mem[0487] = 000;
  font_mem[0488] = 006;
  font_mem[0489] = 000;
  font_mem[0490] = 000;
  font_mem[0491] = 006;
  font_mem[0492] = 024;
  font_mem[0493] = 000;
  font_mem[0494] = 000;
  font_mem[0495] = 000;
  font_mem[0496] = 000;
  font_mem[0497] = 000;
  font_mem[0498] = 000;
  font_mem[0499] = 000;
  font_mem[0500] = 006;
  font_mem[0501] = 000;
  font_mem[0502] = 000;
  font_mem[0503] = 000;
  font_mem[0504] = 000;
  font_mem[0505] = 000;
  font_mem[0506] = 000;
  font_mem[0507] = 012;
  font_mem[0508] = 024;
  font_mem[0509] = 012;
  font_mem[0510] = 115;
  font_mem[0511] = 008;
  font_mem[0512] = 000;
  font_mem[0513] = 000;
  font_mem[0514] = 165;
  font_mem[0515] = 127;
  font_mem[0516] = 127;
  font_mem[0517] = 255;
  font_mem[0518] = 255;
  font_mem[0519] = 000;
  font_mem[0520] = 255;
  font_mem[0521] = 085;
  font_mem[0522] = 069;
  font_mem[0523] = 078;
  font_mem[0524] = 102;
  font_mem[0525] = 054;
  font_mem[0526] = 198;
  font_mem[0527] = 126;
  font_mem[0528] = 124;
  font_mem[0529] = 031;
  font_mem[0530] = 024;
  font_mem[0531] = 102;
  font_mem[0532] = 219;
  font_mem[0533] = 060;
  font_mem[0534] = 000;
  font_mem[0535] = 024;
  font_mem[0536] = 024;
  font_mem[0537] = 024;
  font_mem[0538] = 006;
  font_mem[0539] = 048;
  font_mem[0540] = 003;
  font_mem[0541] = 102;
  font_mem[0542] = 028;
  font_mem[0543] = 062;
  font_mem[0544] = 000;
  font_mem[0545] = 030;
  font_mem[0546] = 036;
  font_mem[0547] = 054;
  font_mem[0548] = 003;
  font_mem[0549] = 051;
  font_mem[0550] = 014;
  font_mem[0551] = 006;
  font_mem[0552] = 006;
  font_mem[0553] = 048;
  font_mem[0554] = 060;
  font_mem[0555] = 024;
  font_mem[0556] = 000;
  font_mem[0557] = 000;
  font_mem[0558] = 000;
  font_mem[0559] = 048;
  font_mem[0560] = 123;
  font_mem[0561] = 012;
  font_mem[0562] = 048;
  font_mem[0563] = 048;
  font_mem[0564] = 054;
  font_mem[0565] = 003;
  font_mem[0566] = 003;
  font_mem[0567] = 096;
  font_mem[0568] = 051;
  font_mem[0569] = 051;
  font_mem[0570] = 028;
  font_mem[0571] = 028;
  font_mem[0572] = 006;
  font_mem[0573] = 126;
  font_mem[0574] = 048;
  font_mem[0575] = 024;
  font_mem[0576] = 123;
  font_mem[0577] = 051;
  font_mem[0578] = 102;
  font_mem[0579] = 003;
  font_mem[0580] = 102;
  font_mem[0581] = 038;
  font_mem[0582] = 038;
  font_mem[0583] = 003;
  font_mem[0584] = 051;
  font_mem[0585] = 012;
  font_mem[0586] = 048;
  font_mem[0587] = 054;
  font_mem[0588] = 006;
  font_mem[0589] = 127;
  font_mem[0590] = 111;
  font_mem[0591] = 099;
  font_mem[0592] = 102;
  font_mem[0593] = 099;
  font_mem[0594] = 102;
  font_mem[0595] = 003;
  font_mem[0596] = 012;
  font_mem[0597] = 051;
  font_mem[0598] = 051;
  font_mem[0599] = 099;
  font_mem[0600] = 030;
  font_mem[0601] = 051;
  font_mem[0602] = 024;
  font_mem[0603] = 012;
  font_mem[0604] = 006;
  font_mem[0605] = 048;
  font_mem[0606] = 000;
  font_mem[0607] = 000;
  font_mem[0608] = 000;
  font_mem[0609] = 030;
  font_mem[0610] = 062;
  font_mem[0611] = 030;
  font_mem[0612] = 062;
  font_mem[0613] = 030;
  font_mem[0614] = 006;
  font_mem[0615] = 110;
  font_mem[0616] = 054;
  font_mem[0617] = 030;
  font_mem[0618] = 060;
  font_mem[0619] = 102;
  font_mem[0620] = 024;
  font_mem[0621] = 063;
  font_mem[0622] = 031;
  font_mem[0623] = 030;
  font_mem[0624] = 059;
  font_mem[0625] = 110;
  font_mem[0626] = 055;
  font_mem[0627] = 030;
  font_mem[0628] = 063;
  font_mem[0629] = 051;
  font_mem[0630] = 051;
  font_mem[0631] = 099;
  font_mem[0632] = 099;
  font_mem[0633] = 102;
  font_mem[0634] = 063;
  font_mem[0635] = 006;
  font_mem[0636] = 024;
  font_mem[0637] = 024;
  font_mem[0638] = 000;
  font_mem[0639] = 028;
  font_mem[0640] = 000;
  font_mem[0641] = 000;
  font_mem[0642] = 129;
  font_mem[0643] = 127;
  font_mem[0644] = 127;
  font_mem[0645] = 231;
  font_mem[0646] = 255;
  font_mem[0647] = 000;
  font_mem[0648] = 000;
  font_mem[0649] = 093;
  font_mem[0650] = 069;
  font_mem[0651] = 031;
  font_mem[0652] = 060;
  font_mem[0653] = 028;
  font_mem[0654] = 198;
  font_mem[0655] = 231;
  font_mem[0656] = 127;
  font_mem[0657] = 127;
  font_mem[0658] = 024;
  font_mem[0659] = 102;
  font_mem[0660] = 222;
  font_mem[0661] = 102;
  font_mem[0662] = 000;
  font_mem[0663] = 024;
  font_mem[0664] = 024;
  font_mem[0665] = 024;
  font_mem[0666] = 127;
  font_mem[0667] = 127;
  font_mem[0668] = 003;
  font_mem[0669] = 255;
  font_mem[0670] = 028;
  font_mem[0671] = 062;
  font_mem[0672] = 000;
  font_mem[0673] = 012;
  font_mem[0674] = 000;
  font_mem[0675] = 054;
  font_mem[0676] = 030;
  font_mem[0677] = 024;
  font_mem[0678] = 095;
  font_mem[0679] = 000;
  font_mem[0680] = 006;
  font_mem[0681] = 048;
  font_mem[0682] = 255;
  font_mem[0683] = 126;
  font_mem[0684] = 000;
  font_mem[0685] = 127;
  font_mem[0686] = 000;
  font_mem[0687] = 024;
  font_mem[0688] = 107;
  font_mem[0689] = 012;
  font_mem[0690] = 024;
  font_mem[0691] = 028;
  font_mem[0692] = 051;
  font_mem[0693] = 031;
  font_mem[0694] = 031;
  font_mem[0695] = 048;
  font_mem[0696] = 030;
  font_mem[0697] = 062;
  font_mem[0698] = 000;
  font_mem[0699] = 000;
  font_mem[0700] = 003;
  font_mem[0701] = 000;
  font_mem[0702] = 096;
  font_mem[0703] = 012;
  font_mem[0704] = 123;
  font_mem[0705] = 051;
  font_mem[0706] = 062;
  font_mem[0707] = 003;
  font_mem[0708] = 102;
  font_mem[0709] = 062;
  font_mem[0710] = 062;
  font_mem[0711] = 003;
  font_mem[0712] = 063;
  font_mem[0713] = 012;
  font_mem[0714] = 048;
  font_mem[0715] = 030;
  font_mem[0716] = 006;
  font_mem[0717] = 107;
  font_mem[0718] = 127;
  font_mem[0719] = 099;
  font_mem[0720] = 062;
  font_mem[0721] = 099;
  font_mem[0722] = 062;
  font_mem[0723] = 014;
  font_mem[0724] = 012;
  font_mem[0725] = 051;
  font_mem[0726] = 051;
  font_mem[0727] = 107;
  font_mem[0728] = 012;
  font_mem[0729] = 030;
  font_mem[0730] = 012;
  font_mem[0731] = 012;
  font_mem[0732] = 012;
  font_mem[0733] = 048;
  font_mem[0734] = 000;
  font_mem[0735] = 000;
  font_mem[0736] = 000;
  font_mem[0737] = 048;
  font_mem[0738] = 102;
  font_mem[0739] = 051;
  font_mem[0740] = 051;
  font_mem[0741] = 051;
  font_mem[0742] = 031;
  font_mem[0743] = 051;
  font_mem[0744] = 110;
  font_mem[0745] = 024;
  font_mem[0746] = 048;
  font_mem[0747] = 054;
  font_mem[0748] = 024;
  font_mem[0749] = 107;
  font_mem[0750] = 051;
  font_mem[0751] = 051;
  font_mem[0752] = 102;
  font_mem[0753] = 051;
  font_mem[0754] = 118;
  font_mem[0755] = 051;
  font_mem[0756] = 006;
  font_mem[0757] = 051;
  font_mem[0758] = 051;
  font_mem[0759] = 099;
  font_mem[0760] = 054;
  font_mem[0761] = 102;
  font_mem[0762] = 049;
  font_mem[0763] = 003;
  font_mem[0764] = 000;
  font_mem[0765] = 048;
  font_mem[0766] = 000;
  font_mem[0767] = 054;
  font_mem[0768] = 000;
  font_mem[0769] = 000;
  font_mem[0770] = 189;
  font_mem[0771] = 127;
  font_mem[0772] = 062;
  font_mem[0773] = 231;
  font_mem[0774] = 126;
  font_mem[0775] = 000;
  font_mem[0776] = 000;
  font_mem[0777] = 077;
  font_mem[0778] = 069;
  font_mem[0779] = 051;
  font_mem[0780] = 024;
  font_mem[0781] = 028;
  font_mem[0782] = 198;
  font_mem[0783] = 231;
  font_mem[0784] = 124;
  font_mem[0785] = 031;
  font_mem[0786] = 024;
  font_mem[0787] = 000;
  font_mem[0788] = 216;
  font_mem[0789] = 102;
  font_mem[0790] = 000;
  font_mem[0791] = 024;
  font_mem[0792] = 024;
  font_mem[0793] = 024;
  font_mem[0794] = 006;
  font_mem[0795] = 048;
  font_mem[0796] = 003;
  font_mem[0797] = 102;
  font_mem[0798] = 062;
  font_mem[0799] = 028;
  font_mem[0800] = 000;
  font_mem[0801] = 012;
  font_mem[0802] = 000;
  font_mem[0803] = 054;
  font_mem[0804] = 048;
  font_mem[0805] = 012;
  font_mem[0806] = 123;
  font_mem[0807] = 000;
  font_mem[0808] = 006;
  font_mem[0809] = 048;
  font_mem[0810] = 060;
  font_mem[0811] = 024;
  font_mem[0812] = 000;
  font_mem[0813] = 000;
  font_mem[0814] = 000;
  font_mem[0815] = 012;
  font_mem[0816] = 111;
  font_mem[0817] = 012;
  font_mem[0818] = 012;
  font_mem[0819] = 048;
  font_mem[0820] = 127;
  font_mem[0821] = 048;
  font_mem[0822] = 051;
  font_mem[0823] = 024;
  font_mem[0824] = 051;
  font_mem[0825] = 024;
  font_mem[0826] = 000;
  font_mem[0827] = 000;
  font_mem[0828] = 006;
  font_mem[0829] = 126;
  font_mem[0830] = 048;
  font_mem[0831] = 012;
  font_mem[0832] = 123;
  font_mem[0833] = 063;
  font_mem[0834] = 102;
  font_mem[0835] = 003;
  font_mem[0836] = 102;
  font_mem[0837] = 038;
  font_mem[0838] = 038;
  font_mem[0839] = 115;
  font_mem[0840] = 051;
  font_mem[0841] = 012;
  font_mem[0842] = 051;
  font_mem[0843] = 054;
  font_mem[0844] = 070;
  font_mem[0845] = 099;
  font_mem[0846] = 123;
  font_mem[0847] = 099;
  font_mem[0848] = 006;
  font_mem[0849] = 115;
  font_mem[0850] = 054;
  font_mem[0851] = 024;
  font_mem[0852] = 012;
  font_mem[0853] = 051;
  font_mem[0854] = 051;
  font_mem[0855] = 107;
  font_mem[0856] = 030;
  font_mem[0857] = 012;
  font_mem[0858] = 006;
  font_mem[0859] = 012;
  font_mem[0860] = 024;
  font_mem[0861] = 048;
  font_mem[0862] = 000;
  font_mem[0863] = 000;
  font_mem[0864] = 000;
  font_mem[0865] = 062;
  font_mem[0866] = 102;
  font_mem[0867] = 003;
  font_mem[0868] = 051;
  font_mem[0869] = 063;
  font_mem[0870] = 006;
  font_mem[0871] = 051;
  font_mem[0872] = 102;
  font_mem[0873] = 024;
  font_mem[0874] = 048;
  font_mem[0875] = 030;
  font_mem[0876] = 024;
  font_mem[0877] = 107;
  font_mem[0878] = 051;
  font_mem[0879] = 051;
  font_mem[0880] = 102;
  font_mem[0881] = 051;
  font_mem[0882] = 110;
  font_mem[0883] = 006;
  font_mem[0884] = 006;
  font_mem[0885] = 051;
  font_mem[0886] = 051;
  font_mem[0887] = 107;
  font_mem[0888] = 028;
  font_mem[0889] = 102;
  font_mem[0890] = 024;
  font_mem[0891] = 006;
  font_mem[0892] = 024;
  font_mem[0893] = 024;
  font_mem[0894] = 000;
  font_mem[0895] = 099;
  font_mem[0896] = 000;
  font_mem[0897] = 000;
  font_mem[0898] = 153;
  font_mem[0899] = 062;
  font_mem[0900] = 028;
  font_mem[0901] = 024;
  font_mem[0902] = 024;
  font_mem[0903] = 000;
  font_mem[0904] = 000;
  font_mem[0905] = 085;
  font_mem[0906] = 093;
  font_mem[0907] = 051;
  font_mem[0908] = 126;
  font_mem[0909] = 054;
  font_mem[0910] = 230;
  font_mem[0911] = 126;
  font_mem[0912] = 112;
  font_mem[0913] = 007;
  font_mem[0914] = 126;
  font_mem[0915] = 000;
  font_mem[0916] = 216;
  font_mem[0917] = 060;
  font_mem[0918] = 127;
  font_mem[0919] = 126;
  font_mem[0920] = 024;
  font_mem[0921] = 126;
  font_mem[0922] = 012;
  font_mem[0923] = 024;
  font_mem[0924] = 127;
  font_mem[0925] = 036;
  font_mem[0926] = 062;
  font_mem[0927] = 028;
  font_mem[0928] = 000;
  font_mem[0929] = 000;
  font_mem[0930] = 000;
  font_mem[0931] = 127;
  font_mem[0932] = 048;
  font_mem[0933] = 006;
  font_mem[0934] = 051;
  font_mem[0935] = 000;
  font_mem[0936] = 012;
  font_mem[0937] = 024;
  font_mem[0938] = 102;
  font_mem[0939] = 024;
  font_mem[0940] = 000;
  font_mem[0941] = 000;
  font_mem[0942] = 000;
  font_mem[0943] = 006;
  font_mem[0944] = 103;
  font_mem[0945] = 012;
  font_mem[0946] = 006;
  font_mem[0947] = 048;
  font_mem[0948] = 048;
  font_mem[0949] = 048;
  font_mem[0950] = 051;
  font_mem[0951] = 012;
  font_mem[0952] = 051;
  font_mem[0953] = 024;
  font_mem[0954] = 028;
  font_mem[0955] = 028;
  font_mem[0956] = 012;
  font_mem[0957] = 000;
  font_mem[0958] = 024;
  font_mem[0959] = 000;
  font_mem[0960] = 003;
  font_mem[0961] = 051;
  font_mem[0962] = 102;
  font_mem[0963] = 099;
  font_mem[0964] = 102;
  font_mem[0965] = 006;
  font_mem[0966] = 006;
  font_mem[0967] = 099;
  font_mem[0968] = 051;
  font_mem[0969] = 012;
  font_mem[0970] = 051;
  font_mem[0971] = 054;
  font_mem[0972] = 102;
  font_mem[0973] = 099;
  font_mem[0974] = 115;
  font_mem[0975] = 099;
  font_mem[0976] = 006;
  font_mem[0977] = 123;
  font_mem[0978] = 102;
  font_mem[0979] = 051;
  font_mem[0980] = 012;
  font_mem[0981] = 051;
  font_mem[0982] = 051;
  font_mem[0983] = 054;
  font_mem[0984] = 051;
  font_mem[0985] = 012;
  font_mem[0986] = 070;
  font_mem[0987] = 012;
  font_mem[0988] = 048;
  font_mem[0989] = 048;
  font_mem[0990] = 000;
  font_mem[0991] = 000;
  font_mem[0992] = 000;
  font_mem[0993] = 051;
  font_mem[0994] = 102;
  font_mem[0995] = 003;
  font_mem[0996] = 051;
  font_mem[0997] = 003;
  font_mem[0998] = 006;
  font_mem[0999] = 051;
  font_mem[1000] = 102;
  font_mem[1001] = 024;
  font_mem[1002] = 048;
  font_mem[1003] = 054;
  font_mem[1004] = 024;
  font_mem[1005] = 107;
  font_mem[1006] = 051;
  font_mem[1007] = 051;
  font_mem[1008] = 102;
  font_mem[1009] = 051;
  font_mem[1010] = 006;
  font_mem[1011] = 024;
  font_mem[1012] = 006;
  font_mem[1013] = 051;
  font_mem[1014] = 051;
  font_mem[1015] = 107;
  font_mem[1016] = 028;
  font_mem[1017] = 102;
  font_mem[1018] = 006;
  font_mem[1019] = 012;
  font_mem[1020] = 024;
  font_mem[1021] = 012;
  font_mem[1022] = 000;
  font_mem[1023] = 099;
  font_mem[1024] = 000;
  font_mem[1025] = 000;
  font_mem[1026] = 195;
  font_mem[1027] = 028;
  font_mem[1028] = 008;
  font_mem[1029] = 024;
  font_mem[1030] = 024;
  font_mem[1031] = 000;
  font_mem[1032] = 000;
  font_mem[1033] = 034;
  font_mem[1034] = 034;
  font_mem[1035] = 051;
  font_mem[1036] = 024;
  font_mem[1037] = 099;
  font_mem[1038] = 231;
  font_mem[1039] = 219;
  font_mem[1040] = 096;
  font_mem[1041] = 003;
  font_mem[1042] = 060;
  font_mem[1043] = 102;
  font_mem[1044] = 216;
  font_mem[1045] = 048;
  font_mem[1046] = 127;
  font_mem[1047] = 060;
  font_mem[1048] = 024;
  font_mem[1049] = 060;
  font_mem[1050] = 000;
  font_mem[1051] = 000;
  font_mem[1052] = 000;
  font_mem[1053] = 000;
  font_mem[1054] = 127;
  font_mem[1055] = 008;
  font_mem[1056] = 000;
  font_mem[1057] = 012;
  font_mem[1058] = 000;
  font_mem[1059] = 054;
  font_mem[1060] = 031;
  font_mem[1061] = 051;
  font_mem[1062] = 059;
  font_mem[1063] = 000;
  font_mem[1064] = 024;
  font_mem[1065] = 012;
  font_mem[1066] = 000;
  font_mem[1067] = 000;
  font_mem[1068] = 028;
  font_mem[1069] = 000;
  font_mem[1070] = 028;
  font_mem[1071] = 003;
  font_mem[1072] = 099;
  font_mem[1073] = 012;
  font_mem[1074] = 051;
  font_mem[1075] = 051;
  font_mem[1076] = 048;
  font_mem[1077] = 051;
  font_mem[1078] = 051;
  font_mem[1079] = 012;
  font_mem[1080] = 051;
  font_mem[1081] = 012;
  font_mem[1082] = 028;
  font_mem[1083] = 028;
  font_mem[1084] = 024;
  font_mem[1085] = 000;
  font_mem[1086] = 012;
  font_mem[1087] = 012;
  font_mem[1088] = 003;
  font_mem[1089] = 051;
  font_mem[1090] = 102;
  font_mem[1091] = 102;
  font_mem[1092] = 054;
  font_mem[1093] = 070;
  font_mem[1094] = 006;
  font_mem[1095] = 102;
  font_mem[1096] = 051;
  font_mem[1097] = 012;
  font_mem[1098] = 051;
  font_mem[1099] = 102;
  font_mem[1100] = 102;
  font_mem[1101] = 099;
  font_mem[1102] = 099;
  font_mem[1103] = 054;
  font_mem[1104] = 006;
  font_mem[1105] = 062;
  font_mem[1106] = 102;
  font_mem[1107] = 051;
  font_mem[1108] = 012;
  font_mem[1109] = 051;
  font_mem[1110] = 030;
  font_mem[1111] = 054;
  font_mem[1112] = 051;
  font_mem[1113] = 012;
  font_mem[1114] = 099;
  font_mem[1115] = 012;
  font_mem[1116] = 096;
  font_mem[1117] = 048;
  font_mem[1118] = 000;
  font_mem[1119] = 000;
  font_mem[1120] = 000;
  font_mem[1121] = 051;
  font_mem[1122] = 102;
  font_mem[1123] = 051;
  font_mem[1124] = 051;
  font_mem[1125] = 051;
  font_mem[1126] = 006;
  font_mem[1127] = 062;
  font_mem[1128] = 102;
  font_mem[1129] = 024;
  font_mem[1130] = 048;
  font_mem[1131] = 102;
  font_mem[1132] = 024;
  font_mem[1133] = 107;
  font_mem[1134] = 051;
  font_mem[1135] = 051;
  font_mem[1136] = 102;
  font_mem[1137] = 051;
  font_mem[1138] = 006;
  font_mem[1139] = 051;
  font_mem[1140] = 054;
  font_mem[1141] = 051;
  font_mem[1142] = 030;
  font_mem[1143] = 054;
  font_mem[1144] = 054;
  font_mem[1145] = 060;
  font_mem[1146] = 035;
  font_mem[1147] = 012;
  font_mem[1148] = 024;
  font_mem[1149] = 012;
  font_mem[1150] = 000;
  font_mem[1151] = 127;
  font_mem[1152] = 000;
  font_mem[1153] = 255;
  font_mem[1154] = 126;
  font_mem[1155] = 008;
  font_mem[1156] = 000;
  font_mem[1157] = 126;
  font_mem[1158] = 126;
  font_mem[1159] = 000;
  font_mem[1160] = 000;
  font_mem[1161] = 028;
  font_mem[1162] = 028;
  font_mem[1163] = 030;
  font_mem[1164] = 024;
  font_mem[1165] = 000;
  font_mem[1166] = 103;
  font_mem[1167] = 024;
  font_mem[1168] = 064;
  font_mem[1169] = 001;
  font_mem[1170] = 024;
  font_mem[1171] = 102;
  font_mem[1172] = 216;
  font_mem[1173] = 099;
  font_mem[1174] = 127;
  font_mem[1175] = 024;
  font_mem[1176] = 024;
  font_mem[1177] = 024;
  font_mem[1178] = 000;
  font_mem[1179] = 000;
  font_mem[1180] = 000;
  font_mem[1181] = 000;
  font_mem[1182] = 127;
  font_mem[1183] = 008;
  font_mem[1184] = 000;
  font_mem[1185] = 012;
  font_mem[1186] = 000;
  font_mem[1187] = 054;
  font_mem[1188] = 012;
  font_mem[1189] = 049;
  font_mem[1190] = 110;
  font_mem[1191] = 000;
  font_mem[1192] = 048;
  font_mem[1193] = 006;
  font_mem[1194] = 000;
  font_mem[1195] = 000;
  font_mem[1196] = 028;
  font_mem[1197] = 000;
  font_mem[1198] = 028;
  font_mem[1199] = 001;
  font_mem[1200] = 062;
  font_mem[1201] = 063;
  font_mem[1202] = 063;
  font_mem[1203] = 030;
  font_mem[1204] = 120;
  font_mem[1205] = 030;
  font_mem[1206] = 030;
  font_mem[1207] = 012;
  font_mem[1208] = 030;
  font_mem[1209] = 014;
  font_mem[1210] = 000;
  font_mem[1211] = 024;
  font_mem[1212] = 048;
  font_mem[1213] = 000;
  font_mem[1214] = 006;
  font_mem[1215] = 012;
  font_mem[1216] = 062;
  font_mem[1217] = 051;
  font_mem[1218] = 063;
  font_mem[1219] = 060;
  font_mem[1220] = 031;
  font_mem[1221] = 127;
  font_mem[1222] = 015;
  font_mem[1223] = 124;
  font_mem[1224] = 051;
  font_mem[1225] = 030;
  font_mem[1226] = 030;
  font_mem[1227] = 103;
  font_mem[1228] = 127;
  font_mem[1229] = 099;
  font_mem[1230] = 099;
  font_mem[1231] = 028;
  font_mem[1232] = 015;
  font_mem[1233] = 048;
  font_mem[1234] = 103;
  font_mem[1235] = 030;
  font_mem[1236] = 030;
  font_mem[1237] = 030;
  font_mem[1238] = 012;
  font_mem[1239] = 054;
  font_mem[1240] = 051;
  font_mem[1241] = 030;
  font_mem[1242] = 127;
  font_mem[1243] = 060;
  font_mem[1244] = 064;
  font_mem[1245] = 060;
  font_mem[1246] = 000;
  font_mem[1247] = 000;
  font_mem[1248] = 000;
  font_mem[1249] = 110;
  font_mem[1250] = 059;
  font_mem[1251] = 030;
  font_mem[1252] = 110;
  font_mem[1253] = 030;
  font_mem[1254] = 015;
  font_mem[1255] = 048;
  font_mem[1256] = 103;
  font_mem[1257] = 126;
  font_mem[1258] = 051;
  font_mem[1259] = 103;
  font_mem[1260] = 126;
  font_mem[1261] = 099;
  font_mem[1262] = 051;
  font_mem[1263] = 030;
  font_mem[1264] = 062;
  font_mem[1265] = 062;
  font_mem[1266] = 015;
  font_mem[1267] = 030;
  font_mem[1268] = 028;
  font_mem[1269] = 110;
  font_mem[1270] = 012;
  font_mem[1271] = 054;
  font_mem[1272] = 099;
  font_mem[1273] = 048;
  font_mem[1274] = 063;
  font_mem[1275] = 056;
  font_mem[1276] = 024;
  font_mem[1277] = 007;
  font_mem[1278] = 000;
  font_mem[1279] = 000;
  font_mem[1280] = 000;
  font_mem[1281] = 000;
  font_mem[1282] = 000;
  font_mem[1283] = 000;
  font_mem[1284] = 000;
  font_mem[1285] = 000;
  font_mem[1286] = 000;
  font_mem[1287] = 000;
  font_mem[1288] = 000;
  font_mem[1289] = 000;
  font_mem[1290] = 000;
  font_mem[1291] = 000;
  font_mem[1292] = 000;
  font_mem[1293] = 000;
  font_mem[1294] = 003;
  font_mem[1295] = 000;
  font_mem[1296] = 000;
  font_mem[1297] = 000;
  font_mem[1298] = 000;
  font_mem[1299] = 000;
  font_mem[1300] = 000;
  font_mem[1301] = 126;
  font_mem[1302] = 000;
  font_mem[1303] = 126;
  font_mem[1304] = 000;
  font_mem[1305] = 000;
  font_mem[1306] = 000;
  font_mem[1307] = 000;
  font_mem[1308] = 000;
  font_mem[1309] = 000;
  font_mem[1310] = 000;
  font_mem[1311] = 000;
  font_mem[1312] = 000;
  font_mem[1313] = 000;
  font_mem[1314] = 000;
  font_mem[1315] = 000;
  font_mem[1316] = 012;
  font_mem[1317] = 000;
  font_mem[1318] = 000;
  font_mem[1319] = 000;
  font_mem[1320] = 000;
  font_mem[1321] = 000;
  font_mem[1322] = 000;
  font_mem[1323] = 000;
  font_mem[1324] = 006;
  font_mem[1325] = 000;
  font_mem[1326] = 000;
  font_mem[1327] = 000;
  font_mem[1328] = 000;
  font_mem[1329] = 000;
  font_mem[1330] = 000;
  font_mem[1331] = 000;
  font_mem[1332] = 000;
  font_mem[1333] = 000;
  font_mem[1334] = 000;
  font_mem[1335] = 000;
  font_mem[1336] = 000;
  font_mem[1337] = 000;
  font_mem[1338] = 000;
  font_mem[1339] = 012;
  font_mem[1340] = 000;
  font_mem[1341] = 000;
  font_mem[1342] = 000;
  font_mem[1343] = 000;
  font_mem[1344] = 000;
  font_mem[1345] = 000;
  font_mem[1346] = 000;
  font_mem[1347] = 000;
  font_mem[1348] = 000;
  font_mem[1349] = 000;
  font_mem[1350] = 000;
  font_mem[1351] = 000;
  font_mem[1352] = 000;
  font_mem[1353] = 000;
  font_mem[1354] = 000;
  font_mem[1355] = 000;
  font_mem[1356] = 000;
  font_mem[1357] = 000;
  font_mem[1358] = 000;
  font_mem[1359] = 000;
  font_mem[1360] = 000;
  font_mem[1361] = 120;
  font_mem[1362] = 000;
  font_mem[1363] = 000;
  font_mem[1364] = 000;
  font_mem[1365] = 000;
  font_mem[1366] = 000;
  font_mem[1367] = 000;
  font_mem[1368] = 000;
  font_mem[1369] = 000;
  font_mem[1370] = 000;
  font_mem[1371] = 000;
  font_mem[1372] = 000;
  font_mem[1373] = 000;
  font_mem[1374] = 000;
  font_mem[1375] = 255;
  font_mem[1376] = 000;
  font_mem[1377] = 000;
  font_mem[1378] = 000;
  font_mem[1379] = 000;
  font_mem[1380] = 000;
  font_mem[1381] = 000;
  font_mem[1382] = 000;
  font_mem[1383] = 051;
  font_mem[1384] = 000;
  font_mem[1385] = 000;
  font_mem[1386] = 051;
  font_mem[1387] = 000;
  font_mem[1388] = 000;
  font_mem[1389] = 000;
  font_mem[1390] = 000;
  font_mem[1391] = 000;
  font_mem[1392] = 006;
  font_mem[1393] = 048;
  font_mem[1394] = 000;
  font_mem[1395] = 000;
  font_mem[1396] = 000;
  font_mem[1397] = 000;
  font_mem[1398] = 000;
  font_mem[1399] = 000;
  font_mem[1400] = 000;
  font_mem[1401] = 024;
  font_mem[1402] = 000;
  font_mem[1403] = 000;
  font_mem[1404] = 000;
  font_mem[1405] = 000;
  font_mem[1406] = 000;
  font_mem[1407] = 000;
  font_mem[1408] = 000;
  font_mem[1409] = 000;
  font_mem[1410] = 000;
  font_mem[1411] = 000;
  font_mem[1412] = 000;
  font_mem[1413] = 000;
  font_mem[1414] = 000;
  font_mem[1415] = 000;
  font_mem[1416] = 000;
  font_mem[1417] = 000;
  font_mem[1418] = 000;
  font_mem[1419] = 000;
  font_mem[1420] = 000;
  font_mem[1421] = 000;
  font_mem[1422] = 000;
  font_mem[1423] = 000;
  font_mem[1424] = 000;
  font_mem[1425] = 000;
  font_mem[1426] = 000;
  font_mem[1427] = 000;
  font_mem[1428] = 000;
  font_mem[1429] = 000;
  font_mem[1430] = 000;
  font_mem[1431] = 000;
  font_mem[1432] = 000;
  font_mem[1433] = 000;
  font_mem[1434] = 000;
  font_mem[1435] = 000;
  font_mem[1436] = 000;
  font_mem[1437] = 000;
  font_mem[1438] = 000;
  font_mem[1439] = 000;
  font_mem[1440] = 000;
  font_mem[1441] = 000;
  font_mem[1442] = 000;
  font_mem[1443] = 000;
  font_mem[1444] = 000;
  font_mem[1445] = 000;
  font_mem[1446] = 000;
  font_mem[1447] = 000;
  font_mem[1448] = 000;
  font_mem[1449] = 000;
  font_mem[1450] = 000;
  font_mem[1451] = 000;
  font_mem[1452] = 000;
  font_mem[1453] = 000;
  font_mem[1454] = 000;
  font_mem[1455] = 000;
  font_mem[1456] = 000;
  font_mem[1457] = 000;
  font_mem[1458] = 000;
  font_mem[1459] = 000;
  font_mem[1460] = 000;
  font_mem[1461] = 000;
  font_mem[1462] = 000;
  font_mem[1463] = 000;
  font_mem[1464] = 000;
  font_mem[1465] = 000;
  font_mem[1466] = 000;
  font_mem[1467] = 000;
  font_mem[1468] = 000;
  font_mem[1469] = 000;
  font_mem[1470] = 000;
  font_mem[1471] = 000;
  font_mem[1472] = 000;
  font_mem[1473] = 000;
  font_mem[1474] = 000;
  font_mem[1475] = 000;
  font_mem[1476] = 000;
  font_mem[1477] = 000;
  font_mem[1478] = 000;
  font_mem[1479] = 000;
  font_mem[1480] = 000;
  font_mem[1481] = 000;
  font_mem[1482] = 000;
  font_mem[1483] = 000;
  font_mem[1484] = 000;
  font_mem[1485] = 000;
  font_mem[1486] = 000;
  font_mem[1487] = 000;
  font_mem[1488] = 000;
  font_mem[1489] = 000;
  font_mem[1490] = 000;
  font_mem[1491] = 000;
  font_mem[1492] = 000;
  font_mem[1493] = 000;
  font_mem[1494] = 000;
  font_mem[1495] = 000;
  font_mem[1496] = 000;
  font_mem[1497] = 000;
  font_mem[1498] = 000;
  font_mem[1499] = 000;
  font_mem[1500] = 000;
  font_mem[1501] = 000;
  font_mem[1502] = 000;
  font_mem[1503] = 000;
  font_mem[1504] = 000;
  font_mem[1505] = 000;
  font_mem[1506] = 000;
  font_mem[1507] = 000;
  font_mem[1508] = 000;
  font_mem[1509] = 000;
  font_mem[1510] = 000;
  font_mem[1511] = 030;
  font_mem[1512] = 000;
  font_mem[1513] = 000;
  font_mem[1514] = 030;
  font_mem[1515] = 000;
  font_mem[1516] = 000;
  font_mem[1517] = 000;
  font_mem[1518] = 000;
  font_mem[1519] = 000;
  font_mem[1520] = 015;
  font_mem[1521] = 120;
  font_mem[1522] = 000;
  font_mem[1523] = 000;
  font_mem[1524] = 000;
  font_mem[1525] = 000;
  font_mem[1526] = 000;
  font_mem[1527] = 000;
  font_mem[1528] = 000;
  font_mem[1529] = 015;
  font_mem[1530] = 000;
  font_mem[1531] = 000;
  font_mem[1532] = 000;
  font_mem[1533] = 000;
  font_mem[1534] = 000;
  font_mem[1535] = 000;
end

always @(posedge CLK or negedge nRST)
  if (!nRST) begin
    rddata <= 8'h0;
    addr_r <= 11'h00;
    rden_r <= 1'b0;
  end else begin
    addr_r <= {char_line,char_addr};
    rden_r <= rden;

    if (rden_r)
      rddata <= font_mem[addr_r];
  end

endmodule
